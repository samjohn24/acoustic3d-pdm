module top();
   bf_time_pcm_tb_mod tb();
   test_program pgm();
endmodule
